------------------------------------------------------------
-- VHDL Top
-- 2015 2 5 19 36 15
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.10.33625
------------------------------------------------------------

------------------------------------------------------------
-- VHDL Top
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity Top Is
  attribute MacroCell : boolean;

End Top;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of Top Is
   Component Kontakter                                       -- ObjectKind=Sheet Symbol|PrimaryId=CONN
   End Component;



Begin
    CONN : Kontakter                                         -- ObjectKind=Sheet Symbol|PrimaryId=CONN
;

End Structure;
------------------------------------------------------------

