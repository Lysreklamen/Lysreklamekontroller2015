------------------------------------------------------------
-- VHDL Kontakter
-- 2015 2 5 19 40 29
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.10.33625
------------------------------------------------------------

------------------------------------------------------------
-- VHDL Kontakter
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity Kontakter Is
  attribute MacroCell : boolean;

End Kontakter;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of Kontakter Is


Begin
End Structure;
------------------------------------------------------------

