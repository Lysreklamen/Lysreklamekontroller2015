------------------------------------------------------------
-- VHDL Bokskort_top
-- 2015 2 5 19 40 29
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 14.3.10.33625
------------------------------------------------------------

------------------------------------------------------------
-- VHDL Bokskort_top
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity Bokskort_top Is
  attribute MacroCell : boolean;

End Bokskort_top;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of Bokskort_top Is
   Component Kontakter                                       -- ObjectKind=Sheet Symbol|PrimaryId=Designator
   End Component;



Begin
    Designator : Kontakter                                   -- ObjectKind=Sheet Symbol|PrimaryId=Designator
;

End Structure;
------------------------------------------------------------

